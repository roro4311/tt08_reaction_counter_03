module tt_um_reaction_timer (
    input wire clk,
    input wire rst_n,
    input wire [7:0] ui_in,
    output wire [7:0] uo_out,
    output wire [7:0] uio_out,
    output wire [7:0] uio_oe,
    input wire [7:0] uio_in,  // Added uio_in port
    input wire ena
);

    wire miso, cs;
    wire [7:0] data_out;

    // SPI driver instance
    spi_driver spi_inst (
        .clk(clk),
        .rst_n(rst_n),
        .miso(miso),
        .cs(cs),
        .data_out(data_out)
    );
 // Instantiate the reaction_timer module
    reaction_timer reaction_timer_inst (
        .clk(clk),
        .rst_n(rst_n),
        .ena(ena),
        .ui_in(ui_in),
        .uo_out(uo_out), // Adjust connections as needed
        .uio_out(uio_out), // Adjust connections as needed
        .uio_oe(uio_oe) // Adjust connections as needed
    );

    // Logic to connect ui_in and handle outputs
    assign uo_out = 8'b0; // Assign outputs as needed

    // Assuming uio_oe is used for controlling tri-state outputs
    assign uio_oe = 8'b11111111; // Example: set all as outputs

    // Connect data_out from SPI driver to uio_out if needed
    assign uio_out = (ena) ? data_out : 8'b0;

    // Debugging
    initial begin
        $monitor("At time %t, ui_in = %h, miso = %b, cs = %b, data_out = %h, uo_out = %h, uio_out = %h, uio_oe = %h", $time, ui_in, miso, cs, data_out, uo_out, uio_out, uio_oe);
    end

    // Additional logic goes here

endmodule
